//                              -*- Mode: Verilog -*-
// Filename        : RTLTopModule.sv
// Description     : RTL top module (DUT).
// Author          : Adrian Fiergolski
// Created On      : Thu Sep 18 10:50:28 2014
// Last Modified By: Adrian Fiergolski
// Last Modified On: Thu Sep 18 10:50:28 2014
// Update Count    : 0
// Status          : Unknown, Use with caution!

module RTLTopModule;
   includeModule incl();
   ipcore ip();
endmodule // RTLTopModule
